package opcodes;

    parameter NOP = 8'h00;
    parameter HLT = 8'hFF;
    
endpackage